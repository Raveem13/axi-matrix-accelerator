module mac (
    input  logic clk,
    input  logic rst,
    input  logic signed [15:0] a,
    input  logic signed [15:0] b,
    input  logic en,
    output logic signed [31:0] y
);
endmodule