module controller_fsm (
    input  logic clk,
    input  logic rst,
    input  logic start,
    output logic done
);
endmodule
