module top (
    input logic clk,
    input logic rst
);
endmodule
